module core(
    input logic clk,
    input logic rst_n
);

endmodule