module cpu_top(
    input logic clk,
    input logic rst_n
);

endmodule